package sharedpkg ;
bit test_finished ;

int error_cntr = 0  ;
int correct_cntr = 0; 
    
endpackage